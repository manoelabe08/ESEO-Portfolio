
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.Virgule_pkg.all;

entity SegmentDisplayController is
    generic(
        -- Declarations
    );
    port(
        -- Declarations
    );
end SegmentDisplayController;

architecture Behavioral of SegmentDisplayController is
    -- Declarations
begin
    -- Concurrent statements
end Behavioral;
