
architecture Simple of EventDetector is
    -- Declarations
    signal src_reg : std_logic_vector(0 to 1) := "00";
begin
    -- Concurrent statements
end Simple;
