../../c/Loader/Loader_pkg.vhd