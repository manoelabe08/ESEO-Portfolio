
architecture Debouncer of EventDetector is
    -- Declarations
begin
    -- Concurrent statements
end Debouncer;
