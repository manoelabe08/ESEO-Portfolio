
library ieee;
use ieee.std_logic_1164.all;

entity Pomodoro is
   -- Ports
end Pomodoro;

architecture Structural of Pomodoro is
   -- Declarations.
begin
   -- Concurrent statements.
end Structural;
